`define CSR_REGS    32'h1000_0000
